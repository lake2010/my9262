library verilog;
use verilog.vl_types.all;
entity Verilog_First_vlg_tst is
end Verilog_First_vlg_tst;
