library verilog;
use verilog.vl_types.all;
entity Verilog_First_vlg_check_tst is
    port(
        LED1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Verilog_First_vlg_check_tst;
